library IEEE;
use IEEE.std_logic_1164.all;


entity clo is

	port(
	i_rs : in std_logic_vector(31 downto 0);	--Data being Read in from rs
	o_rd : out std_logic_vector(31 downto 0));	--Amount of 1s

end clo;


architecture dataflow of clo is 

begin


	o_rd <= "00000000000000000000000000100000" when i_rs(31 downto 0) ="11111111111111111111111111111111"	else--32
			"00000000000000000000000000011111" when i_rs(31 downto 1) ="1111111111111111111111111111111"	else--31
			"00000000000000000000000000011110" when i_rs(31 downto 2) ="111111111111111111111111111111"	else--30
			"00000000000000000000000000011101" when i_rs(31 downto 3) ="11111111111111111111111111111"	else--29
			"00000000000000000000000000011100" when i_rs(31 downto 4) ="1111111111111111111111111111"	else--28
			"00000000000000000000000000011011" when i_rs(31 downto 5) ="111111111111111111111111111"	else--27
			"00000000000000000000000000011010" when i_rs(31 downto 6) ="11111111111111111111111111"	else--26
			"00000000000000000000000000011001" when i_rs(31 downto 7) ="1111111111111111111111111"	else--25
			"00000000000000000000000000011000" when i_rs(31 downto 8) ="111111111111111111111111"	else--24
			"00000000000000000000000000010111" when i_rs(31 downto 9) ="11111111111111111111111"	else--23
			"00000000000000000000000000010110" when i_rs(31 downto 10)="1111111111111111111111"	else--22
			"00000000000000000000000000010101" when i_rs(31 downto 11)="111111111111111111111"	else--21
			"00000000000000000000000000010100" when i_rs(31 downto 12)="11111111111111111111"	else--20
			"00000000000000000000000000010011" when i_rs(31 downto 13)="1111111111111111111"	else--19
			"00000000000000000000000000010010" when i_rs(31 downto 14)="111111111111111111"					else--18
			"00000000000000000000000000010001" when i_rs(31 downto 15)="11111111111111111"					else--17
			"00000000000000000000000000010000" when i_rs(31 downto 16)="1111111111111111"					else--16
			"00000000000000000000000000001111" when i_rs(31 downto 17)="111111111111111"					else--15
			"00000000000000000000000000001110" when i_rs(31 downto 18)="11111111111111"						else--18
			"00000000000000000000000000001101" when i_rs(31 downto 19)="1111111111111"						else--13
			"00000000000000000000000000001100" when i_rs(31 downto 20)="111111111111"						else--12
			"00000000000000000000000000001011" when i_rs(31 downto 21)="11111111111"						else--11
			"00000000000000000000000000001010" when i_rs(31 downto 22)="1111111111"							else--10
			"00000000000000000000000000001001" when i_rs(31 downto 23)="111111111"							else--9
			"00000000000000000000000000001000" when i_rs(31 downto 24)="11111111"							else--8
			"00000000000000000000000000000111" when i_rs(31 downto 25)="1111111"							else--7
			"00000000000000000000000000000110" when i_rs(31 downto 26)="111111"							else--6
			"00000000000000000000000000000101" when i_rs(31 downto 27)="11111"							else--5
			"00000000000000000000000000000100" when i_rs(31 downto 28)="1111"							else--4
			"00000000000000000000000000000011" when i_rs(31 downto 29)="111"							else--3
			"00000000000000000000000000000010" when i_rs(31 downto 30)="11"							else--2
			"00000000000000000000000000000001" when i_rs(31)		  ='1'							else--1

			"00000000000000000000000000000000";


end dataflow;
